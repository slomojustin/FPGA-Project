module control_block_fetch (
    input [31:0] pc,
    output bios_ena
);

assign bios_ena = 1'b1;

endmodule